------------------------------------------------
-- Project:	Sudoku - Game
------------------------------------------------
-- Entity:	rom_lbl
-- Date:		31.05.2016
-- Description:
-- 	ROM with Bit-Matrix of Labels
------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_lbl is
	generic(
		ROM_WIDTH	: natural := 128;	-- count of columns
		ROM_DEPTH	: natural := 32;	-- count of rows
		ADR_WIDTH	: natural := 9		-- address width -> label(4-bit) + line(5-bit)
	);
	port(
		rom_adr_i	: in	std_logic_vector(ADR_WIDTH - 1 downto 0);
		rom_dat_o	: out std_logic_vector(ROM_WIDTH - 1 downto 0)
	);
end rom_lbl;

architecture rtl of rom_lbl is
	
	subtype rom_row_t is std_logic_vector(0 to ROM_WIDTH - 1);
	type rom_mem_t is array(0 to ROM_DEPTH - 1) of rom_row_t;
	
	constant rom_lbl_start : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "00000000000000000000000000000000111111110000000011000000000000000000000000000000000000000011000000000000000000000000000000000000",
		 9 => "00000000000000000000000000000001110000010000000011000000000000000000000000000000000000000011000000000000000000000000000000000000",
		10 => "00000000000000000000000000000011000000000000000011000000000000000000000000000000000000000011000000000000000000000000000000000000",
		11 => "00000000000000000000000000000011000000000000000011000000000000000000000000000000000000000011000000000000000000000000000000000000",
		12 => "00000000000000000000000000000011000000000000111111111110000001111110000000011001111000111111111110000000000000000000000000000000",
		13 => "00000000000000000000000000000011000000000000111111111110000011111111100000011011111100111111111110000000000000000000000000000000",
		14 => "00000000000000000000000000000001110000000000000011000000000011000001100000011110000100000011000000000000000000000000000000000000",
		15 => "00000000000000000000000000000001111110000000000011000000000000000000110000011100000000000011000000000000000000000000000000000000",
		16 => "00000000000000000000000000000000011111100000000011000000000000000000110000011000000000000011000000000000000000000000000000000000",
		17 => "00000000000000000000000000000000000001110000000011000000000000111111110000011000000000000011000000000000000000000000000000000000",
		18 => "00000000000000000000000000000000000000111000000011000000000011111111110000011000000000000011000000000000000000000000000000000000",
		19 => "00000000000000000000000000000000000000011000000011000000000111000000110000011000000000000011000000000000000000000000000000000000",
		20 => "00000000000000000000000000000000000000011000000011000000000110000000110000011000000000000011000000000000000000000000000000000000",
		21 => "00000000000000000000000000000000000000011000000011000000000110000001110000011000000000000011000000000000000000000000000000000000",
		22 => "00000000000000000000000000000011000001110000000011100000000111000011110000011000000000000011100000000000000000000000000000000000",
		23 => "00000000000000000000000000000011111111110000000001111110000011111110110000011000000000000001111110000000000000000000000000000000",
		24 => "00000000000000000000000000000001111111000000000000111110000001111100110000011000000000000000111110000000000000000000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		
	constant rom_lbl_restart : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000011100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "00000000011100000011000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000011000000000000000",
		 9 => "00000000011110000011000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000011000000000000000",
		10 => "00000000011110000011000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000011000000000000000",
		11 => "00000000011011000011000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000011000000000000000",
		12 => "00000000011011000011000000011111000000110000000110000011111110000111111111110000001111110000000011001111000111111111110000000000",
		13 => "00000000011011000011000000111111110000110000000110000111111111000111111111110000011111111100000011011111100111111111110000000000",
		14 => "00000000011001100011000001110000110000110000000110001110000001000000011000000000011000001100000011110000100000011000000000000000",
		15 => "00000000011001100011000001100000011000110000000110001100000000000000011000000000000000000110000011100000000000011000000000000000",
		16 => "00000000011000110011000011000000011000110000000110001110000000000000011000000000000000000110000011000000000000011000000000000000",
		17 => "00000000011000110011000011111111111000110000000110000111111000000000011000000000000111111110000011000000000000011000000000000000",
		18 => "00000000011000011011000011111111111000110000000110000011111111000000011000000000011111111110000011000000000000011000000000000000",
		19 => "00000000011000011011000011000000000000110000000110000000001111100000011000000000111000000110000011000000000000011000000000000000",
		20 => "00000000011000011011000011000000000000110000000110000000000001100000011000000000110000000110000011000000000000011000000000000000",
		21 => "00000000011000001111000001100000000000110000001110000000000001100000011000000000110000001110000011000000000000011000000000000000",
		22 => "00000000011000001111000001110000010000111000011110001100000011100000011100000000111000011110000011000000000000011100000000000000",
		23 => "00000000011000000111000000111111110000011111110110001111111111000000001111110000011111110110000011000000000000001111110000000000",
		24 => "00000000011000000111000000011111100000001111100110000011111100000000000111110000001111100110000011000000000000000111110000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");


	constant rom_lbl_exit : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000000000001111111000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000",
		 8 => "00000000000000001111111110000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000",
		 9 => "00000000000000001100000110000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000",
		10 => "00000000000000001100000011000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000",
		11 => "00000000000000001100000011000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000",
		12 => "00000000000000001100000011000000001111100000000011111000000110011111000000001111001100000011111000000110011111000000000000000000",
		13 => "00000000000000001100000011000000011111111000000111111110000110111111100000011111111100000111111110000110111111100000000000000000",
		14 => "00000000000000001100000110000000111000011000001110000110000111100001110000111000111100001110000110000111100001110000000000000000",
		15 => "00000000000000001111111100000000110000001100001100000011000111000000110001110000011100001100000011000111000000110000000000000000",
		16 => "00000000000000001111111110000001100000001100011000000011000110000000110001100000001100011000000011000110000000110000000000000000",
		17 => "00000000000000001100000111000001111111111100011111111111000110000000110001100000001100011111111111000110000000110000000000000000",
		18 => "00000000000000001100000001100001111111111100011111111111000110000000110001100000001100011111111111000110000000110000000000000000",
		19 => "00000000000000001100000001100001100000000000011000000000000110000000110001100000001100011000000000000110000000110000000000000000",
		20 => "00000000000000001100000001100001100000000000011000000000000110000000110001100000001100011000000000000110000000110000000000000000",
		21 => "00000000000000001100000001100000110000000000001100000000000110000000110001110000011100001100000000000110000000110000000000000000",
		22 => "00000000000000001100000011100000111000001000001110000010000110000000110000111000111100001110000010000110000000110000000000000000",
		23 => "00000000000000001111111111000000011111111000000111111110000110000000110000011111111100000111111110000110000000110000000000000000",
		24 => "00000000000000001111111100000000001111110000000011111100000110000000110000001111001100000011111100000110000000110000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

	constant rom_lbl_difficulty : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000011000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000011000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000",
		 7 => "00000000000000000000000000011000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000",
		 8 => "00000000000000000000000000011000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000",
		 9 => "00000000000000000000000000011000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000",
		10 => "00000000000000000000000000011000000000000000011111000000110000000110000001111100000000011000000000000000000000000000000000000000",
		11 => "00000000000000000000000000011000000000000000111111110000111000001110000011111111000000011000000000000011100000000000000000000000",
		12 => "00000000000000000000000000011000000000000001110000110000011000001100000111000011000000011000000000000011100000000000000000000000",
		13 => "00000000000000000000000000011000000000000001100000011000011000001100000110000001100000011000000000000011100000000000000000000000",
		14 => "00000000000000000000000000011000000000000011000000011000011100011100001100000001100000011000000000000011100000000000000000000000",
		15 => "00000000000000000000000000011000000000000011111111111000001100011000001111111111100000011000000000000000000000000000000000000000",
		16 => "00000000000000000000000000011000000000000011111111111000001100011000001111111111100000011000000000000000000000000000000000000000",
		17 => "00000000000000000000000000011000000000000011000000000000001110111000001100000000000000011000000000000000000000000000000000000000",
		18 => "00000000000000000000000000011000000000000011000000000000000110110000001100000000000000011000000000000000000000000000000000000000",
		19 => "00000000000000000000000000011000000000000001100000000000000110110000000110000000000000011000000000000011100000000000000000000000",
		20 => "00000000000000000000000000011000000000000001110000010000000111110000000111000001000000011100000000000011100000000000000000000000",
		21 => "00000000000000000000000000011111111111000000111111110000000011100000000011111111000000001111110000000011100000000000000000000000",
		22 => "00000000000000000000000000011111111111000000011111100000000011100000000001111110000000000111110000000011100000000000000000000000",
		23 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		24 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		

	constant rom_lbl_easy : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000000000000000000110000000000000000000000000000000110000000000000000000000110000000000000000000000000000000000000000000000",
		 8 => "00000000000000000000000110000000000000000000000000000000110000000000000000000000110000000000000001100000000000000000000000000000",
		 9 => "00000000000000000000000110000000000000000000000000000000110000000000000000000000110000000000000001100000000000000000000000000000",
		10 => "00000000000000000000000110000000000000000000000000000000000000000000000000000000110000000000000001100000000000000001111000000000",
		11 => "00000000000000000000000110000000000000000000000000000000000000000000000000000000110000000000000001100000000000000000111100000000",
		12 => "00000000000000000000000110000000000000000111110000000111110000000000001111100000110011111000011111111111000000000000011110000000",
		13 => "00000000000000000000000110000000000000001111111100000111110000000000111111110000110111111100011111111111000000000000001111000000",
		14 => "00000000000000000000000110000000000000011100001100000000110000000001110000010000111100001110000001100000000000000000000111100000",
		15 => "00000000000000000000000110000000000000011000000110000000110000000001100000000000111000000110000001100000000000000000000011110000",
		16 => "00000000000000000000000110000000000000110000000110000000110000000011000000000000110000000110000001100000000000000000000001111000",
		17 => "00000000000000000000000110000000000000111111111110000000110000000011000000000000110000000110000001100000000000000000000011110000",
		18 => "00000000000000000000000110000000000000111111111110000000110000000011000000000000110000000110000001100000000000000000000111100000",
		19 => "00000000000000000000000110000000000000110000000000000000110000000011000000000000110000000110000001100000000000000000001111000000",
		20 => "00000000000000000000000110000000000000110000000000000000110000000011000000000000110000000110000001100000000000000000011110000000",
		21 => "00000000000000000000000110000000000000011000000000000000110000000001100000000000110000000110000001100000000000000000111100000000",
		22 => "00000000000000000000000110000000000000011100000100000000110000000001110000010000110000000110000001110000000000000001111000000000",
		23 => "00000000000000000000000111111111110000001111111100001111111111000000111111110000110000000110000000111111000000000000000000000000",
		24 => "00000000000000000000000111111111110000000111111000001111111111000000001111100000110000000110000000011111000000000000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

	constant rom_lbl_medium : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000000000000000000111000000111000000011000000000000000000000000000000000000000000000000011111100000000000000000000000000000",
		 8 => "00000000000000000000000111000000111000000011000000000001100000000000011000000000000000000000011111100000000000000000000000000000",
		 9 => "00000000000000000000000111100001111000000011000000000001100000000000011000000000000000000000000001100000000000000000000000000000",
		10 => "00000000011110000000000111100001111000000000000000000001100000000000011000000000000000000000000001100000000000000001111000000000",
		11 => "00000000111100000000000110100001011000000000000000000001100000000000011000000000000000000000000001100000000000000000111100000000",
		12 => "00000001111000000000000110110011011000011111000000011111111111000111111111110000000111110000000001100000000000000000011110000000",
		13 => "00000011110000000000000110110011011000011111000000011111111111000111111111110000001111111100000001100000000000000000001111000000",
		14 => "00000111100000000000000110010010011000000011000000000001100000000000011000000000011100001100000001100000000000000000000111100000",
		15 => "00001111000000000000000110011110011000000011000000000001100000000000011000000000011000000110000001100000000000000000000011110000",
		16 => "00011110000000000000000110011110011000000011000000000001100000000000011000000000110000000110000001100000000000000000000001111000",
		17 => "00001111000000000000000110001100011000000011000000000001100000000000011000000000111111111110000001100000000000000000000011110000",
		18 => "00000111100000000000000110001100011000000011000000000001100000000000011000000000111111111110000001100000000000000000000111100000",
		19 => "00000011110000000000000110000000011000000011000000000001100000000000011000000000110000000000000001100000000000000000001111000000",
		20 => "00000001111000000000000110000000011000000011000000000001100000000000011000000000110000000000000001100000000000000000011110000000",
		21 => "00000000111100000000000110000000011000000011000000000001100000000000011000000000011000000000000001100000000000000000111100000000",
		22 => "00000000011110000000000110000000011000000011000000000001110000000000011100000000011100000100000001110000000000000001111000000000",
		23 => "00000000000000000000000110000000011000111111111100000000111111000000001111110000001111111100000000111111000000000000000000000000",
		24 => "00000000000000000000000110000000011000111111111100000000011111000000000111110000000111111000000000011111000000000000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

	constant rom_lbl_hard : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000000000000000000000111111000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "00000000000000000000000001111111100000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000",
		 9 => "00000000000000000000000011100000100000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000",
		10 => "00000000011110000000000110000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000",
		11 => "00000000111100000000000110000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000",
		12 => "00000001111000000000000110000000000000000011111000001100111110001100000000001100000111110000000011001111000000000000000000000000",
		13 => "00000011110000000000000110000000000000001111111100001101111111001100000000001100001111111100000011011111100000000000000000000000",
		14 => "00000111100000000000000011100000000000011100000100001111000011100110000000011000011100001100000011110000100000000000000000000000",
		15 => "00001111000000000000000011111100000000011000000000001110000001100110000000011000011000000110000011100000000000000000000000000000",
		16 => "00011110000000000000000000111111000000110000000000001100000001100110001100011000110000000110000011000000000000000000000000000000",
		17 => "00001111000000000000000000000011100000110000000000001100000001100110001100011000111111111110000011000000000000000000000000000000",
		18 => "00000111100000000000000000000001110000110000000000001100000001100111011110111000111111111110000011000000000000000000000000000000",
		19 => "00000011110000000000000000000000110000110000000000001100000001100011011110110000110000000000000011000000000000000000000000000000",
		20 => "00000001111000000000000000000000110000110000000000001100000001100011010010110000110000000000000011000000000000000000000000000000",
		21 => "00000000111100000000000000000000110000011000000000001100000001100011110011110000011000000000000011000000000000000000000000000000",
		22 => "00000000011110000000000110000011100000011100000100001100000001100011110011110000011100000100000011000000000000000000000000000000",
		23 => "00000000000000000000000111111111100000001111111100001100000001100001100001100000001111111100000011000000000000000000000000000000",
		24 => "00000000000000000000000011111110000000000011111000001100000001100001100001100000000111111000000011000000000000000000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
	
	constant rom_lbl_sudoku : rom_mem_t := (
		 0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 9 => "00000000000000000000000000000001111000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000",
		10 => "00000000000000000000000000000010000100000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000",
		11 => "00000000000000000000000000000100000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000",
		12 => "00000000000000000000000000000100000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000",
		13 => "00000000000000000000000000000100000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000",
		14 => "00000000000000000000000000000010000000000000000000000000001000000000000001000000000000000000000000000000000000000000000000000000",
		15 => "00000000000000000000000000000001111000001000000100000111101000001111000001000001100010000001000000000000000000000000000000000000",
		16 => "00000000000000000000000000000000000100001000000100001000011000010000100001000110000010000001000000000000000000000000000000000000",
		17 => "00000000000000000000000000000000000010001000000100010000001000100000010001011000000010000001000000000000000000000000000000000000",
		18 => "00000000000000000000000000000000000010001000000100010000001000100000010001100000000010000001000000000000000000000000000000000000",
		19 => "00000000000000000000000000000000000010001000000100010000001000100000010001011000000010000001000000000000000000000000000000000000",
		20 => "00000000000000000000000000000010000100000100001100001000011000010000100001000110000001000011000000000000000000000000000000000000",
		21 => "00000000000000000000000000000001111000000011110100000111101000001111000001000001100000111101000000000000000000000000000000000000",
		22 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		23 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		24 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		25 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		28 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		29 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		30 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		31 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		
	signal bit_dat	: std_logic_vector(0 to ROM_WIDTH - 1);
	signal lbl_adr	: std_logic_vector(3 downto 0);
	signal bit_adr	: std_logic_vector(4 downto 0);
	
begin
	
	lbl_adr <= rom_adr_i(8 downto 5);
	bit_adr <= rom_adr_i(4 downto 0);
	
	process(lbl_adr, bit_adr, bit_dat)
	begin
		case lbl_adr is
			when "0001" => bit_dat <= rom_lbl_start(to_integer(unsigned(bit_adr)));
			when "0010" => bit_dat <= rom_lbl_restart(to_integer(unsigned(bit_adr)));
			when "0011" => bit_dat <= rom_lbl_exit(to_integer(unsigned(bit_adr)));
			when "0100" => bit_dat <= rom_lbl_difficulty(to_integer(unsigned(bit_adr)));
			when "0101" => bit_dat <= rom_lbl_easy(to_integer(unsigned(bit_adr)));
			when "0110" => bit_dat <= rom_lbl_medium(to_integer(unsigned(bit_adr)));
			when "0111" => bit_dat <= rom_lbl_hard(to_integer(unsigned(bit_adr)));
			when "1000" => bit_dat <= rom_lbl_sudoku(to_integer(unsigned(bit_adr)));
			when others => bit_dat <= (others => '0');
		end case;
		
		rom_dat_o <= bit_dat;
	end process;
end rtl;
------------------------------------------------
-- Project:	Sudoku - Game
------------------------------------------------
-- Entity:	rom_mem
-- Date:		07.05.2016
-- Description:
-- 	ROM with Bit-Matrix of Numbers
------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_mem is
	generic(
		ROM_WIDTH	: natural := 32;	-- count of columns
		ROM_DEPTH	: natural := 32;	-- count of rows
		ADR_WIDTH	: natural := 9		-- address width -> number(4-bit) + line(5-bit)
	);
	port(
		rom_adr_i	: in	std_logic_vector(ADR_WIDTH - 1 downto 0);
		rom_dat_o	: out std_logic_vector(ROM_WIDTH - 1 downto 0)
	);
end rom_mem;

architecture rtl of rom_mem is
	
	subtype rom_row_t is std_logic_vector(0 to ROM_WIDTH - 1);
	type rom_mem_t is array(0 to ROM_DEPTH - 1) of rom_row_t;
	
	constant rom_mdl_1 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000001111110000000000000",
		 6 => "00000000000111111110000000000000",
		 7 => "00000000000111111110000000000000",
		 8 => "00000000000111001110000000000000",
		 9 => "00000000000000001110000000000000",
		10 => "00000000000000001110000000000000",
		11 => "00000000000000001110000000000000",
		12 => "00000000000000001110000000000000",
		13 => "00000000000000001110000000000000",
		14 => "00000000000000001110000000000000",
		15 => "00000000000000001110000000000000",
		16 => "00000000000000001110000000000000",
		17 => "00000000000000001110000000000000",
		18 => "00000000000000001110000000000000",
		19 => "00000000000000001110000000000000",
		20 => "00000000000000001110000000000000",
		21 => "00000000000000001110000000000000",
		22 => "00000000000000001110000000000000",
		23 => "00000000000000001110000000000000",
		24 => "00000000000111111111111100000000",
		25 => "00000000000111111111111100000000",
		26 => "00000000000111111111111100000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_2 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000011111111000000000000",
		 6 => "00000000001111111111110000000000",
		 7 => "00000000001111111111111000000000",
		 8 => "00000000001100000001111000000000",
		 9 => "00000000000000000000111100000000",
		10 => "00000000000000000000011100000000",
		11 => "00000000000000000000011100000000",
		12 => "00000000000000000000011100000000",
		13 => "00000000000000000000011100000000",
		14 => "00000000000000000000111100000000",
		15 => "00000000000000000001111000000000",
		16 => "00000000000000000011110000000000",
		17 => "00000000000000000111110000000000",
		18 => "00000000000000001111000000000000",
		19 => "00000000000000011110000000000000",
		20 => "00000000000000111100000000000000",
		21 => "00000000000001111000000000000000",
		22 => "00000000000011110000000000000000",
		23 => "00000000000111000000000000000000",
		24 => "00000000001111111111111100000000",
		25 => "00000000001111111111111100000000",
		26 => "00000000001111111111111100000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_3 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000011111100000000000000",
		 6 => "00000000001111111111000000000000",
		 7 => "00000000001111111111100000000000",
		 8 => "00000000001100000111110000000000",
		 9 => "00000000000000000001110000000000",
		10 => "00000000000000000001110000000000",
		11 => "00000000000000000001110000000000",
		12 => "00000000000000000001110000000000",
		13 => "00000000000000000111100000000000",
		14 => "00000000000001111111000000000000",
		15 => "00000000000001111110000000000000",
		16 => "00000000000001111111100000000000",
		17 => "00000000000000000011110000000000",
		18 => "00000000000000000001110000000000",
		19 => "00000000000000000000111000000000",
		20 => "00000000000000000000111000000000",
		21 => "00000000000000000000111000000000",
		22 => "00000000000000000001111000000000",
		23 => "00000000011000000011110000000000",
		24 => "00000000011111111111110000000000",
		25 => "00000000011111111111100000000000",
		26 => "00000000000111111110000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_4 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000000000111100000000000",
		 6 => "00000000000000000111100000000000",
		 7 => "00000000000000001111100000000000",
		 8 => "00000000000000011111100000000000",
		 9 => "00000000000000011011100000000000",
		10 => "00000000000000111011100000000000",
		11 => "00000000000000110011100000000000",
		12 => "00000000000001100011100000000000",
		13 => "00000000000011100011100000000000",
		14 => "00000000000011000011100000000000",
		15 => "00000000000111000011100000000000",
		16 => "00000000000110000011100000000000",
		17 => "00000000001110000011100000000000",
		18 => "00000000011100000011100000000000",
		19 => "00000000011111111111111100000000",
		20 => "00000000011111111111111100000000",
		21 => "00000000011111111111111100000000",
		22 => "00000000000000000011100000000000",
		23 => "00000000000000000011100000000000",
		24 => "00000000000000000011100000000000",
		25 => "00000000000000000011100000000000",
		26 => "00000000000000000011100000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_5 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000001111111111100000000000",
		 6 => "00000000001111111111100000000000",
		 7 => "00000000001111111111100000000000",
		 8 => "00000000001110000000000000000000",
		 9 => "00000000001110000000000000000000",
		10 => "00000000001110000000000000000000",
		11 => "00000000001110000000000000000000",
		12 => "00000000001110000000000000000000",
		13 => "00000000001111111110000000000000",
		14 => "00000000001111111111000000000000",
		15 => "00000000001111111111110000000000",
		16 => "00000000001000000111110000000000",
		17 => "00000000000000000001111000000000",
		18 => "00000000000000000000111000000000",
		19 => "00000000000000000000111000000000",
		20 => "00000000000000000000111000000000",
		21 => "00000000000000000000111000000000",
		22 => "00000000000000000001111000000000",
		23 => "00000000011000000011110000000000",
		24 => "00000000011111111111100000000000",
		25 => "00000000011111111111000000000000",
		26 => "00000000000111111100000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_6 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000000111111000000000000",
		 6 => "00000000000011111111100000000000",
		 7 => "00000000000111111111100000000000",
		 8 => "00000000000111100000100000000000",
		 9 => "00000000001111000000000000000000",
		10 => "00000000001110000000000000000000",
		11 => "00000000011110000000000000000000",
		12 => "00000000011100000000000000000000",
		13 => "00000000011100011110000000000000",
		14 => "00000000011101111111100000000000",
		15 => "00000000011101111111110000000000",
		16 => "00000000011111000011110000000000",
		17 => "00000000011110000001111000000000",
		18 => "00000000011100000000111000000000",
		19 => "00000000011100000000111000000000",
		20 => "00000000011100000000111000000000",
		21 => "00000000001100000000111000000000",
		22 => "00000000001110000001111000000000",
		23 => "00000000001111000011110000000000",
		24 => "00000000000111111111110000000000",
		25 => "00000000000011111111100000000000",
		26 => "00000000000001111110000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_7 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000011111111111111000000000",
		 6 => "00000000011111111111111000000000",
		 7 => "00000000011111111111111000000000",
		 8 => "00000000000000000001110000000000",
		 9 => "00000000000000000001110000000000",
		10 => "00000000000000000011100000000000",
		11 => "00000000000000000011100000000000",
		12 => "00000000000000000111100000000000",
		13 => "00000000000000000111000000000000",
		14 => "00000000000000000111000000000000",
		15 => "00000000000000001111000000000000",
		16 => "00000000000000001110000000000000",
		17 => "00000000000000001110000000000000",
		18 => "00000000000000011100000000000000",
		19 => "00000000000000011100000000000000",
		20 => "00000000000000111100000000000000",
		21 => "00000000000000111000000000000000",
		22 => "00000000000000111000000000000000",
		23 => "00000000000001111000000000000000",
		24 => "00000000000001110000000000000000",
		25 => "00000000000001110000000000000000",
		26 => "00000000000011100000000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_8 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000001111110000000000000",
		 6 => "00000000000011111111000000000000",
		 7 => "00000000000111111111100000000000",
		 8 => "00000000001111000011110000000000",
		 9 => "00000000001110000001110000000000",
		10 => "00000000001110000001110000000000",
		11 => "00000000001110000001110000000000",
		12 => "00000000001110000001110000000000",
		13 => "00000000000111000011100000000000",
		14 => "00000000000011111111000000000000",
		15 => "00000000000001111110000000000000",
		16 => "00000000000111111111100000000000",
		17 => "00000000001111000011110000000000",
		18 => "00000000001110000001110000000000",
		19 => "00000000011100000000111000000000",
		20 => "00000000011100000000111000000000",
		21 => "00000000011100000000111000000000",
		22 => "00000000011110000001111000000000",
		23 => "00000000011111000011110000000000",
		24 => "00000000001111111111110000000000",
		25 => "00000000000111111111100000000000",
		26 => "00000000000001111110000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	constant rom_mdl_9 : rom_mem_t := (
		 0 => "00000000000000000000000000000000",
		 1 => "00000000000000000000000000000000",
		 2 => "00000000000000000000000000000000",
		 3 => "00000000000000000000000000000000",
		 4 => "00000000000000000000000000000000",
		 5 => "00000000000011111100000000000000",
		 6 => "00000000001111111110000000000000",
		 7 => "00000000011111111111000000000000",
		 8 => "00000000011110000111100000000000",
		 9 => "00000000111100000011100000000000",
		10 => "00000000111000000001100000000000",
		11 => "00000000111000000001110000000000",
		12 => "00000000111000000001110000000000",
		13 => "00000000111000000001110000000000",
		14 => "00000000111100000011110000000000",
		15 => "00000000011110000111110000000000",
		16 => "00000000011111111101110000000000",
		17 => "00000000001111111101110000000000",
		18 => "00000000000011110001110000000000",
		19 => "00000000000000000001110000000000",
		20 => "00000000000000000011110000000000",
		21 => "00000000000000000011100000000000",
		22 => "00000000000000000111100000000000",
		23 => "00000000001000001111000000000000",
		24 => "00000000001111111111000000000000",
		25 => "00000000001111111110000000000000",
		26 => "00000000000111111000000000000000",
		27 => "00000000000000000000000000000000",
		28 => "00000000000000000000000000000000",
		29 => "00000000000000000000000000000000",
		30 => "00000000000000000000000000000000",
		31 => "00000000000000000000000000000000");
	
	signal bit_dat	: std_logic_vector(0 to ROM_WIDTH - 1);
	signal num_adr	: std_logic_vector(3 downto 0);
	signal bit_adr	: std_logic_vector(4 downto 0);
	
begin
	
	num_adr <= rom_adr_i(8 downto 5);
	bit_adr <= rom_adr_i(4 downto 0);
	
	process(num_adr, bit_adr, bit_dat)
	begin
		case num_adr is
			when "0001" => bit_dat <= rom_mdl_1(to_integer(unsigned(bit_adr)));
			when "0010" => bit_dat <= rom_mdl_2(to_integer(unsigned(bit_adr)));
			when "0011" => bit_dat <= rom_mdl_3(to_integer(unsigned(bit_adr)));
			when "0100" => bit_dat <= rom_mdl_4(to_integer(unsigned(bit_adr)));
			when "0101" => bit_dat <= rom_mdl_5(to_integer(unsigned(bit_adr)));
			when "0110" => bit_dat <= rom_mdl_6(to_integer(unsigned(bit_adr)));
			when "0111" => bit_dat <= rom_mdl_7(to_integer(unsigned(bit_adr)));
			when "1000" => bit_dat <= rom_mdl_8(to_integer(unsigned(bit_adr)));
			when "1001" => bit_dat <= rom_mdl_9(to_integer(unsigned(bit_adr)));
			when others => bit_dat <= (others => '0');
		end case;
		
		rom_dat_o <= bit_dat;
	end process;
end rtl;
------------------------------------------------
-- Project:	Sudoku - Game
------------------------------------------------
-- Entity:	rom_lbl_header
-- Date:		03.06.2016
-- Description:
-- 	ROM with Bit-Matrix of Header-Labels
------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_lbl_header is
	generic(
		ROM_WIDTH	: natural := 256;	-- count of columns
		ROM_DEPTH	: natural := 64;	-- count of rows
		ADR_WIDTH	: natural := 10	-- address width -> label(4-bit) + line(6-bit)
	);
	port(
		rom_adr_i	: in	std_logic_vector(ADR_WIDTH - 1 downto 0);
		rom_dat_o	: out std_logic_vector(ROM_WIDTH - 1 downto 0)
	);
end rom_lbl_header;

architecture rtl of rom_lbl_header is
	
	subtype rom_row_t is std_logic_vector(0 to ROM_WIDTH - 1);
	type rom_mem_t is array(0 to ROM_DEPTH - 1) of rom_row_t;
	
	constant rom_lbl_sudoku : rom_mem_t := (
		 0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000",
		 9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000",
		10 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000",
		11 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000",
		12 => "0000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000",
		13 => "0000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000",
		14 => "0000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		15 => "0000000000000000000000000000000000000000000000000000000000000000110000011111100000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		16 => "0000000000000000000000000000000000000000000000000000000000000011100000001111100000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		17 => "0000000000000000000000000000000000000000000000000000000000000011000000001111100000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		18 => "0000000000000000000000000000000000000000000000000000000000000110000000000111000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		19 => "0000000000000000000000000000000000000000000000000000000000001110000000000100000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		20 => "0000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		21 => "0000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		22 => "0000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		23 => "0000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000111100000000001111100000000000000000000000000000000000000000000000000000000000000000000",
		24 => "0000000000000000000000000000000000000000000000000000000000111100000000000000000000000000110000000000001000000000000000000011111111000000000000000000000111110000000000001111100000000011111110000000000110000000000001000000000000000000000000000000000000000000",
		25 => "0000000000000000000000000000000000000000000000000000000000111110000000000000000000000011110000000000110000000000000000001111111111000000000000000000111111111000000000001111000000000111111100000000011110000000000110000000000000000000000000000000000000000000",
		26 => "0000000000000000000000000000000000000000000000000000000000111110000000000000000000001111110000000011110000000000000000111111111111000000000000000011111111111100000000001111000000001111111000000001111110000000011110000000000000000000000000000000000000000000",
		27 => "0000000000000000000000000000000000000000000000000000000000111111000000000000000000011111100000000011110000000000000001110001111111000000000000000111000011111110000000001111000000011000111000000011111100000000011110000000000000000000000000000000000000000000",
		28 => "0000000000000000000000000000000000000000000000000000000000111111100000000000000001111111100000000011110000000000000111000000011110000000000000011110000001111110000000011111000000110000000000001111111100000000011110000000000000000000000000000000000000000000",
		29 => "0000000000000000000000000000000000000000000000000000000000011111110000000000000011000111100000000111100000000000001110000000011110000000000000111100000001111110000000011110000011100000000000011000111100000000111100000000000000000000000000000000000000000000",
		30 => "0000000000000000000000000000000000000000000000000000000000011111111000000000000000000111100000000111100000000000011110000000011110000000000001111000000000111110000000011110000111000000000000000000111100000000111100000000000000000000000000000000000000000000",
		31 => "0000000000000000000000000000000000000000000000000000000000001111111100000000000000000111000000000111100000000000011100000000111110000000000011110000000000111110000000011110001110000000000000000000111000000000111100000000000000000000000000000000000000000000",
		32 => "0000000000000000000000000000000000000000000000000000000000000111111110000000000000001111000000000111000000000000111100000000111100000000000111100000000000111110000000011110011100000000000000000001111000000000111000000000000000000000000000000000000000000000",
		33 => "0000000000000000000000000000000000000000000000000000000000000011111111100000000000001111000000001111000000000001111000000000111100000000000111100000000000111110000000111110111000000000000000000001111000000001111000000000000000000000000000000000000000000000",
		34 => "0000000000000000000000000000000000000000000000000000000000000001111111100000000000001111000000001111000000000001111000000000111100000000001111100000000000111100000000111101111000000000000000000001111000000001111000000000000000000000000000000000000000000000",
		35 => "0000000000000000000000000000000000000000000000000000000000000000111111110000000000001111000000001111000000000001111000000000111100000000001111000000000000111100000000111111111000000000000000000001111000000001111000000000000000000000000000000000000000000000",
		36 => "0000000000000000000000000000000000000000000000000000000000000000011111111000000000011110000000001110000000000011110000000001111100000000001111000000000000111100000000111111111100000000000000000011110000000001110000000000000000000000000000000000000000000000",
		37 => "0000000000000000000000000000000000000000000000000000000000000000001111111000000000011110000000011110000000000011110000000001111000000000011111000000000001111100000001111101111100000000000000000011110000000011110000000000000000000000000000000000000000000000",
		38 => "0000000000000000000000000000000000000000000000000000000000000000000111111000000000011110000000011110000000000011110000000001111000000000011110000000000001111000000001111000111110000000000000000011110000000011110000000000000000000000000000000000000000000000",
		39 => "0000000000000000000000000000000000000000000000000000000000000000000111111000000000011110000000011110000000000111110000000001111000000000011110000000000001111000000001111000111110000000000000000011110000000011110000000000000000000000000000000000000000000000",
		40 => "0000000000000000000000000000000000000000000000000000000000000000000011111000000000111100000000011110000000000111100000000011111000000000111110000000000011110000000001111000111111000000000000000111100000000011110000000000000000000000000000000000000000000000",
		41 => "0000000000000000000000000000000000000000000000000000000000000000000011111000000000111100000000111100000000000111100000000011111000000000111110000000000011110000000001111000011111000000000000000111100000000111100000000000000000000000000000000000000000000000",
		42 => "0000000000000000000000000000000000000000000000000000000000000000000011110000000000111100000001111100000000000111100000000011110000000000111110000000000111100000000011110000011111100000000000000111100000001111100000000000000000000000000000000000000000000000",
		43 => "0000000000000000000000000000000000000000000000001000000000000000000011110000000000111100000111111100000011001111100000001111110000000100111110000000000111100000000011110000001111100000000000000111100000111111100000011000000000000000000000000000000000000000",
		44 => "0000000000000000000000000000000000000000000000011000000000000000000011100000000001111100001110111100001110001111100000011111110000011100111110000000001111000000000011110000001111100000000000001111100001110111100001110000000000000000000000000000000000000000",
		45 => "0000000000000000000000000000000000000000000000011000000000000000000111100000000001111100111100111100111000001111100001111111110000110000111111000000001110000000000011110000000111110000000000001111100111100111100111000000000000000000000000000000000000000000",
		46 => "0000000000000000000000000000000000000000000000011100000000000000000111000000000001111111110001111111110000001111110011100111110011100000111111000000011100000000000111110000000111110000000000001111111110001111111110000000000000000000000000000000000000000000",
		47 => "0000000000000000000000000000000000000000000000111100000000000000001110000000000001111111100001111111100000001111111110000111111110000000011111100001110000000000000111100000000111111000000000001111111100001111111100000000000000000000000000000000000000000000",
		48 => "0000000000000000000000000000000000000000000000111110000000000000001100000000000001111110000001111110000000001111111100000111111000000000011111111111100000000000000111100000000011111000000000001111110000001111110000000000000000000000000000000000000000000000",
		49 => "0000000000000000000000000000000000000000000001111111000000000000011100000000000001111100000001111000000000000111110000000111110000000000001111111110000000000000000111000000000011111100000000001111100000001111000000000000000000000000000000000000000000000000",
		50 => "0000000000000000000000000000000000000000000001111111100000000001110000000000000000110000000001110000000000000011000000000111000000000000000111110000000000000000000000000000000001111100000000000110000000001110000000000000000000000000000000000000000000000000",
		51 => "0000000000000000000000000000000000000000000000111111111000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000",
		52 => "0000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000",
		53 => "0000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000",
		54 => "0000000000000000000000000000000000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000100000000000000000000000000000000000000000000000000000000000",
		55 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000001100000000000000000000000000000000000000000000000000000000000",
		56 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000011110000000000000000000000000000000000000000000000000000000000",
		57 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000111110000000000000000000000000000000000000000000000000000000000",
		58 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000",
		59 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000",
		60 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		61 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		62 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		63 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		
	constant rom_lbl_credits : rom_mem_t := (
		 0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		10 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		11 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		12 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		13 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		14 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		15 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		16 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		17 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		18 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		19 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		20 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		21 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000",
		22 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
		23 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000110000010000000000000000000000000000000000000000000000000000000000000001111000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
		24 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000001110011100000100000110000000000000000000000000000000000000000001110000000000000000010011000000000000000000000110000000000000000000000000000000000000000000000000000000000000",
		25 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000010000011100001100000110000000000000000000000001000000000000000100110000000000000000100001000001000000000000000110000000000000000000000000000000000000000000000000000000000000",
		26 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101100001100000100000000000000000000000011000000000000001000100000010000000001100000000011000000000000000100000000000000000000000000000000000000000000000000000000000000",
		27 => "0000000000000000000000000000000000000000000000000011000000000000000000000000000000110000101100001000001100000000000000000000000011000000000000011101000000010000000001100000000011000000000000001100000000000000000000000000000000000000000000000000000000000000",
		28 => "0000000000000000000000000000000000000000000111110011000000111000001000110000000000110001001100001000001100110000001100000101100010000000000000001110111111100000000001100000000010000000011000001100000001111000001000110000000000000000000000000000000000000000",
		29 => "0000000000000000000000000000000000000000001000100011000010011100111011100000000000000010001000011000001101111000110110011111111111110000000001001000100110000000000001110000001111110001101101111111000110011000111011100000000000000000000000000000000000000000",
		30 => "0000000000000000000000000000000000000000001001000010000100001100011100100000000000000100001000011000001100011001100100001100000110000000000010100001000100000000000000111000000110000011001000001000001100011000011100100000000000000000000000000000000000000000",
		31 => "0000000000000000000000000000000000000000000011000010001100001100011001100000000000000111111000011000011000011001001000001000000110000000000011000000001100000000000000011100000110000010010000001000001000011000011001100000000000000000000000000000000000000000",
		32 => "0000000000000000000000000000000000000000000010000100011000001000110001100000000000001111111000010000011000010011110000001000000100000000000110000000001000000000000000001110000100000111100000011000001000010000110001100000000000000000000000000000000000000000",
		33 => "0000000000000000000000000000000000000000000110000100011000011000110001000000000000011000011000110000011000110011000000011000000100000000000110000000010000000000000000000110000100000110000000011000011000110000110001000000000000000000000000000000000000000000",
		34 => "0000000000000000000000000000000000000000000110001000011000010000110001000000000000100000011000110010010000100011000000011000001100100000000110000000100000000000000000000100001100100110000000010000011001110100110001000000000000000000000000000000000000000000",
		35 => "0000000000000000000000000000000000000000000111110000011100100000100011001000000111000000011000111000011011000011101000010000001111000000000011100011000000000000010000000100001111000111010000010000011110111000100011001000000000000000000000000000000000000000",
		36 => "0000000000000000000000000000000000000000000011000000001110000001100011100000001110000000011100110000111100000001110000010000000100000000000001111100000000000000110000001000000100000011100000110000011000100001100011100000000000000000000000000000000000000000",
		37 => "0000000000000000000000000000000000000000000000000000000000000001000011000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000111100010000000000000000000000100000000000000001000011000000000000000000000000000000000000000000",
		38 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
		39 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
		40 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
		41 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
		42 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000",
		43 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		44 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		45 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		46 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		47 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		48 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		49 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		50 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		51 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		52 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		53 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		54 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		55 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		56 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		57 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		58 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		59 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		60 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		61 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		62 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		63 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		
	constant rom_lbl_game_won : rom_mem_t := (
		 0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "0000000000000001100000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "0000111000000111100000000000000000000111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "0000111110011111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "0000111111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "0000011111111111000000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "0000011111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "0000011111111111000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 9 => "0000011111111111100000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		10 => "0000111111111111110000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		11 => "0000111111111111111100000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		12 => "0001111111111111111110000000000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		13 => "0011111111111111111110000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		14 => "0111111111111111100000000000000111100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		15 => "0000000111111100000000000000000111100000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		16 => "0000000011111100000000000000000111100000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		17 => "0000000001111100000000000000001111100000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		18 => "0000000000111000001111000000001111000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		19 => "0000000000111000011111100000001111000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		20 => "0000000000010000011111100000001111000000000000000001111111111111000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		21 => "0000000000000000111111100000001110000000000000000000111111111110000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		22 => "0000000000000000111111100000001110000000000000000000011111111100000000000000000000000000111000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		23 => "0000000000000000111111110000001110000000000000110000011111111100000000000000000000000001100000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		24 => "0000000000000000011111110000001100000000000001111000011111111100000000000000000000000011000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		25 => "0000000000000000011111110000001100000000000011111000011111111100000000000000000000000110000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "0000000000000000001111111000001100000000000111110000011100011100000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "0000000000000000000111111000001100000000001111110000010000000100000000000000000000011100000000000000000000000001110000000000000000000000000001110000000001111000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000",
		28 => "0000000000000000000111111000001100000000011111110000000000000000000000000000000000011000000000000000000000000111111000000000000000000000000001110000000111111100000001100000011100000001100000011100000000111111000000011000000111000000000000000000000000000000",
		29 => "0000000000000000000111111000001100000000111111111000000000000000000000000000000000111000000000000000000000001100111000001111111100000110000001110000001100011110000011100000111100000011100000111100000001100111000000111000001111000000000000000000000000000000",
		30 => "0000000000000000000011111000001100000000111111111000000000000000000000000000000000110000000000000000000000011000111000011111111100001110000001110000110000011110001111100011111000001111100011111000000011000111000011111000111110000000000000000000000000000000",
		31 => "0000000000000000000011111100001000000001111111110000000000000000000000000000000001110000000000000000000000110000111000011000011000001110000001110001100000001110010011001110111000010011001110111000000110000111000100110011101110000000000000000000000000000000",
		32 => "0000000000000000000001111100001000000011111111100000000000000000000000000000000001110000000111111111000001110000110000110000110000001100000001100011100000001110000011111000111000000011111000111000001110000110000000111110001110000000000000000000000000000000",
		33 => "0000000000000000000001111100000000000011111111000000000000000000000000000000000001100000001111111110000001100001100000100000100000011100000011100011000000001110000011100000111000000011100000111000001100001100000000111000001110000000000000000000000000000000",
		34 => "0000000000000000000001111100000000000111111110000000000000000000000000000000000011100000000000011100000011100011000000100001100000011100000011000111000000001100000111000000110000000111000000110000011100011000000001110000001100000000000000000000000000000000",
		35 => "0000000000100000000000111100000000000111111100000000000000000000000000000000000011100000000000011100000011100110000000000011000000011000000011000111000000001100000111000000110000000111000000110000011100110000000001110000001100000000000000000000000000000000",
		36 => "0000000001100000000000111110000000001111111000000000000000000000000000000000000011100000000000011000000011011000000000000011000000111000000110000110000000011100000111000001110000000111000001110000011011000000000001110000011100000000000000000000000000000000",
		37 => "0000111111100000000000111110000000001111111000000000000000000000000000000000000011100000000000111000000111110000000000000111000000111000000110001110000000011000000110000001110000000110000001110000111110000000000001100000011100000000000000000000000000000000",
		38 => "0000111111100000000000011110000000011111110000000000000000000000000000000000000011100000000000111000000111000000000000000110000001110000001100001110000000011000001110000001100000001110000001100000111000000000000011100000011000000000000000000000000000000000",
		39 => "0000011111111000000000011110000000011111100000000000000000000000000000000000000011100000000000111000000111000000001000000110000001110000001000001110000000110000001110000001100000001110000001100000111000000001000011100000011000000000000000000000000000000000",
		40 => "0000011111111100000000011110000000011111100000000000000000000000000000000000000011110000000001110000000111000000011000001110000011110000010000001110000000110000001110000001100011001110000001100011111000000011000011100000011000110000000000000000000000000000",
		41 => "0000011111111000000000011110000000111111000000000000000000000000000000000000000001111000000011110000000111000000110000001110000101110000100000001111000001100000001100000011111100001100000011111100111000000110000011000000111111000000000000000000000000000000",
		42 => "0000011111100000000000001110000000111111000000000000000000000000000000000000000001111100001101110000000111100011000000001110011001111001000000001111000010000000011100000011111000011100000011111000111100011000000111000000111110000000000000000000000000000000",
		43 => "0000111111100000010000001110000000111110000000000000000000000000000000000000000000111111110001110000000011111110000000001111110001111110000000000111111100000000011100000011100000011100000011100000011111110000000111000000111000000000000000000000000000000000",
		44 => "0000000001100000111000001110000000111110000000000000000000000000000000000000000000011111000001100000000001111000000000000111000000111000000000000011100000000000000000000010000000000000000010000000001111000000000000000000100000000000000000000000000000000000",
		45 => "0000000000100001111000001111000001111100000000000000000000110000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		46 => "0000000000000001111100000111000001111100000000000000000001110000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		47 => "0000000000000001111100000111000001111000000000000000011111111000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		48 => "0000000000000000111110000111000001111000000000001000001111111110000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		49 => "0000000000000000011110000111000011110000000001111100000111111111000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		50 => "0000000000000000001111000111000011110000000111111100000111111100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		51 => "0000000000000000001111000011000011110000001111111100000111111000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		52 => "0000000000000000000111000011000011100000011111111000001111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		53 => "0000000000000000000111100011000011100000111111000000001100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		54 => "0000000000000000000011100011000011100001111100000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		55 => "0000000000000000000001100011000011000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		56 => "0000000000000000000001100001000011000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		57 => "0000000000000000000001110001000011000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		58 => "0000000000000000000000110001000011001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		59 => "0000000000000000000000110001000010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		60 => "0000000000000000000000010001000010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		61 => "0000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		62 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		63 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		
	constant rom_lbl_game_lost : rom_mem_t := (
		 0 => "0000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 1 => "0000111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 2 => "0001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 3 => "0011111100000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 4 => "0011111000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 5 => "0011110000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 6 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 7 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 8 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		 9 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		10 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		11 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		12 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		13 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		14 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		15 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		16 => "0111100000000000001100000010000000000001000000110000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		17 => "0111100000000000011110000111000000000011100001111000000000000111100000000000000000000000000000000000000000000000000001111000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		18 => "0111100000000000111111001111100000000111110011111100000000000111100000000000000000000000000000000000000000000000000001111000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		19 => "0111100000000000011111111111000000000011111111111000000000000111100000000000000000000000000000000000000000000000000000111000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		20 => "0111100000000000001111111110000000000001111111110000000000000111100000000000000000000000000000000000000000000000000000111000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		21 => "0111100000000000000111111100000000000000111111100000000000000111100000000000000000000000000000000000111111100000000000111000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		22 => "0111100000000000000011111100000000000000111111000000000000000111100000000000000000000000000000000111101111000000000000110000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		23 => "0111100000000000000111111110000000000001111111100000000000000111100000000000000000000000000000001100000111000000000000110000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		24 => "0111100000000000001111111111000000000011111111110000000000000111100000000000000000000000000000011000001111000000000001100000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		25 => "0111100000000000011111111111100000000111111111111000000000000111100000000000000000000000000000110000001110000000000001100000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		26 => "0111100000000000011110001111100000000111110001111000000000000111100000000000000000000000000000110000001110000000000011000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		27 => "0111100000000000001100000111000000000011100000110000000000000111100000000000000000000000000001110000001110000000000110000000001110000000001000011000111000000000000111100000000010000110000000111000000000000000000000000000000000000000000000000000000000000000",
		28 => "0111100000000000000000000010000000000001000000000000000000000111100000000000000000000000000001110000001110000000000100000000111111000000111001111000110000000000011111110000001110011110000011111100000001100000011100000000000000000000000000000000000000000000",
		29 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000001110000001110000000001100000001100111000011111111111001110000000000110001111000111111111110000110011100000011100000111100000000000000000000000000000000000000000000",
		30 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000001111000001110000000011000000011000111001100111100010001110000000011000001111011001111000100001100011100001111100011111000000000000000000000000000000000000000000000",
		31 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000001110000011110000000110000000110000111000000111000000001110000000110000000111000001110000000011000011100010011001110111000000000000000000000000000000000000000000000",
		32 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011100000001100000001110000110000000110000000001100000001110000000111000001100000000111000011000000011111000111000000000000000000000000000000000000000000000",
		33 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011100000001000000001100001100000001110000000011100000001100000000111000011100000000110000110000000011100000111000000000000000000000000000000000000000000000",
		34 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011100000110000000011100011000000001110000000011100000011100000000110000011100000001110001100000000111000000110000000000000000000000000000000000000000000000",
		35 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011100001100000000011100110000000001110000000011100000011100000000110000011100000001110011000000000111000000110000000000000000000000000000000000000000000000",
		36 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011100011000000000011011000000000001100000000011000000011000000001110000011000000001101100000000000111000001110000000000000000000000000000000000000000000000",
		37 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000011100110000000000111110000000000011100000000011000000111000000001100000111000000011111000000000000110000001110000000000000000000000000000000000000000000000",
		38 => "0111100000000000000000000000011111111110000000000000000000000111100000000000000000000000000000000000111001100000000000111000000000000011100000000111000000111000000001100000111000000011100000000000001110000001100000000000000000000000000000000000000000000000",
		39 => "0111100000000000000000000111111111111111110000000000000000000111100000000000000000000000000000000000111011000000000000111000000001000011100000000111000000111000000011000000111000000011100000000100001110000001100000000000000000000000000000000000000000000000",
		40 => "0111100000000000000000111111111111111111111110000000000000000111100000000000000000000000000000000000111110000000000000111000000011000111000000000111000110111000000011000001110000000011100000001100001110000001100011000000000000000000000000000000000000000000",
		41 => "0111100000000000000011111111111111111111111111100000000000000111100000000000000000000000000000000000111100000000000000111000000110000111000000000111001000111100000110000001110000000011100000011000001100000011111100000000000000000000000000000000000000000000",
		42 => "0111100000000000001111111111100000000011111111110000000000000111100000000000000000000000000000000000111000000000000000111100011000000111000000000111110000111100001000000001110000000011110001100000011100000011111000000000000000000000000000000000000000000000",
		43 => "0111100000000000011111111000000000000000001111111000000000000111100000000000000000000000000000000000111000000000000000011111110000000000000000000111100000011111110000000000000000000001111111000000011100000011100000000000000000000000000000000000000000000000",
		44 => "0111100000000000001111100000000000000000000011111000000000000111100000000000000000000000000000000000000000000000000000001111000000000000000000000110000000001110000000000000000000000000111100000000000000000010000000000000000000000000000000000000000000000000",
		45 => "0111100000000000000110000000000000000000000001110000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		46 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		47 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		48 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		49 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		50 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		51 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		52 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		53 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		54 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		55 => "0111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		56 => "0011110000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		57 => "0011111000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		58 => "0011111100000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		59 => "0001111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		60 => "0000111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		61 => "0000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		62 => "0000000011111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
		63 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
		
	signal bit_dat	: std_logic_vector(0 to ROM_WIDTH - 1);
	signal lbl_adr	: std_logic_vector(3 downto 0);
	signal bit_adr	: std_logic_vector(5 downto 0);
	
begin
	
	lbl_adr <= rom_adr_i(9 downto 6);
	bit_adr <= rom_adr_i(5 downto 0);
	
	process(lbl_adr, bit_adr, bit_dat)
	begin
		case lbl_adr is
			when "0001" => bit_dat <= rom_lbl_sudoku(to_integer(unsigned(bit_adr)));
			when "0010" => bit_dat <= rom_lbl_credits(to_integer(unsigned(bit_adr)));
			when "0011" => bit_dat <= rom_lbl_game_won(to_integer(unsigned(bit_adr)));
			when "0100" => bit_dat <= rom_lbl_game_lost(to_integer(unsigned(bit_adr)));
			when others => bit_dat <= (others => '0');
		end case;
		
		rom_dat_o <= bit_dat;
	end process;
end rtl;
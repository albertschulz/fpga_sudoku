------------------------------------------------
-- Project:	Sudoku - Game
------------------------------------------------
-- Entity:	rom_tmr
-- Date:		07.05.2016
-- Description:
-- 	ROM with Bit-Matrix of Numbers for Timer
------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_tmr is
	generic(
		ROM_WIDTH	: natural := 24;	-- count of columns
		ROM_DEPTH	: natural := 32;	-- count of rows
		ADR_WIDTH	: natural := 9		-- address width -> number(4-bit) + line(5-bit)
	);
	port(
		rom_adr_i	: in	std_logic_vector(ADR_WIDTH - 1 downto 0);
		rom_dat_o	: out std_logic_vector(ROM_WIDTH - 1 downto 0)
	);
end rom_tmr;

architecture rtl of rom_tmr is
	
	subtype rom_row_t is std_logic_vector(0 to ROM_WIDTH - 1);
	type rom_mem_t is array(0 to ROM_DEPTH - 1) of rom_row_t;
	
	constant rom_mdl_0 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000000111111000000000",
		 6 => "000000001111111100000000",
		 7 => "000000011111111110000000",
		 8 => "000000111100001111000000",
		 9 => "000000111000000111000000",
		10 => "000001110000000011100000",
		11 => "000001110000000011100000",
		12 => "000001110000000011100000",
		13 => "000001110000000011100000",
		14 => "000001110000000011100000",
		15 => "000001110000000011100000",
		16 => "000001110000000011100000",
		17 => "000001110000000011100000",
		18 => "000001110000000011100000",
		19 => "000001110000000011100000",
		20 => "000001110000000011100000",
		21 => "000001110000000011100000",
		22 => "000001111000000111100000",
		23 => "000001111100001111000000",
		24 => "000000111111111111000000",
		25 => "000000011111111110000000",
		26 => "000000000111111000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
		
	constant rom_mdl_1 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000000111111000000000",
		 6 => "000000011111111000000000",
		 7 => "000000011111111000000000",
		 8 => "000000011100111000000000",
		 9 => "000000000000111000000000",
		10 => "000000000000111000000000",
		11 => "000000000000111000000000",
		12 => "000000000000111000000000",
		13 => "000000000000111000000000",
		14 => "000000000000111000000000",
		15 => "000000000000111000000000",
		16 => "000000000000111000000000",
		17 => "000000000000111000000000",
		18 => "000000000000111000000000",
		19 => "000000000000111000000000",
		20 => "000000000000111000000000",
		21 => "000000000000111000000000",
		22 => "000000000000111000000000",
		23 => "000000000000111000000000",
		24 => "000000011111111111110000",
		25 => "000000011111111111110000",
		26 => "000000011111111111110000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_2 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000011111111000000000",
		 6 => "000001111111111110000000",
		 7 => "000001111111111111000000",
		 8 => "000001100000001111000000",
		 9 => "000000000000000111100000",
		10 => "000000000000000011100000",
		11 => "000000000000000011100000",
		12 => "000000000000000011100000",
		13 => "000000000000000011100000",
		14 => "000000000000000111100000",
		15 => "000000000000001111000000",
		16 => "000000000000011110000000",
		17 => "000000000000111100000000",
		18 => "000000000001111000000000",
		19 => "000000000011110000000000",
		20 => "000000000111100000000000",
		21 => "000000001111000000000000",
		22 => "000000011110000000000000",
		23 => "000000111000000000000000",
		24 => "000001111111111111100000",
		25 => "000001111111111111100000",
		26 => "000001111111111111100000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_3 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000001111110000000000",
		 6 => "000000111111111100000000",
		 7 => "000000111111111110000000",
		 8 => "000000110000011111000000",
		 9 => "000000000000000111000000",
		10 => "000000000000000111000000",
		11 => "000000000000000111000000",
		12 => "000000000000000111000000",
		13 => "000000000000011110000000",
		14 => "000000000111111100000000",
		15 => "000000000111111000000000",
		16 => "000000000111111110000000",
		17 => "000000000000001111000000",
		18 => "000000000000000111000000",
		19 => "000000000000000011100000",
		20 => "000000000000000011100000",
		21 => "000000000000000011100000",
		22 => "000000000000000111100000",
		23 => "000001100000001111000000",
		24 => "000001111111111111000000",
		25 => "000001111111111110000000",
		26 => "000000011111111000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_4 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000000000011110000000",
		 6 => "000000000000011110000000",
		 7 => "000000000000111110000000",
		 8 => "000000000001111110000000",
		 9 => "000000000001101110000000",
		10 => "000000000011101110000000",
		11 => "000000000011001110000000",
		12 => "000000000110001110000000",
		13 => "000000001110001110000000",
		14 => "000000001100001110000000",
		15 => "000000011100001110000000",
		16 => "000000011000001110000000",
		17 => "000000111000001110000000",
		18 => "000001110000001110000000",
		19 => "000001111111111111110000",
		20 => "000001111111111111110000",
		21 => "000001111111111111110000",
		22 => "000000000000001110000000",
		23 => "000000000000001110000000",
		24 => "000000000000001110000000",
		25 => "000000000000001110000000",
		26 => "000000000000001110000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_5 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000111111111110000000",
		 6 => "000000111111111110000000",
		 7 => "000000111111111110000000",
		 8 => "000000111000000000000000",
		 9 => "000000111000000000000000",
		10 => "000000111000000000000000",
		11 => "000000111000000000000000",
		12 => "000000111000000000000000",
		13 => "000000111111111000000000",
		14 => "000000111111111100000000",
		15 => "000000111111111111000000",
		16 => "000000100000011111000000",
		17 => "000000000000000111100000",
		18 => "000000000000000011100000",
		19 => "000000000000000011100000",
		20 => "000000000000000011100000",
		21 => "000000000000000011100000",
		22 => "000000000000000111100000",
		23 => "000001100000001111000000",
		24 => "000001111111111110000000",
		25 => "000001111111111100000000",
		26 => "000000011111110000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_6 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000000011111100000000",
		 6 => "000000001111111110000000",
		 7 => "000000011111111110000000",
		 8 => "000000011110000010000000",
		 9 => "000000111100000000000000",
		10 => "000000111000000000000000",
		11 => "000001111000000000000000",
		12 => "000001110000000000000000",
		13 => "000001110001111000000000",
		14 => "000001110111111110000000",
		15 => "000001110111111111000000",
		16 => "000001111100001111000000",
		17 => "000001111000000111100000",
		18 => "000001110000000011100000",
		19 => "000001110000000011100000",
		20 => "000001110000000011100000",
		21 => "000000110000000011100000",
		22 => "000000111000000111100000",
		23 => "000000111100001111000000",
		24 => "000000011111111111000000",
		25 => "000000001111111110000000",
		26 => "000000000111111000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_7 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000001111111111111100000",
		 6 => "000001111111111111100000",
		 7 => "000001111111111111100000",
		 8 => "000000000000000111000000",
		 9 => "000000000000000111000000",
		10 => "000000000000001110000000",
		11 => "000000000000001110000000",
		12 => "000000000000011110000000",
		13 => "000000000000011100000000",
		14 => "000000000000011100000000",
		15 => "000000000000111100000000",
		16 => "000000000000111000000000",
		17 => "000000000000111000000000",
		18 => "000000000001110000000000",
		19 => "000000000001110000000000",
		20 => "000000000011110000000000",
		21 => "000000000011100000000000",
		22 => "000000000011100000000000",
		23 => "000000000111100000000000",
		24 => "000000000111000000000000",
		25 => "000000000111000000000000",
		26 => "000000000000000000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_8 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000000111111000000000",
		 6 => "000000001111111100000000",
		 7 => "000000011111111110000000",
		 8 => "000000111100001111000000",
		 9 => "000000111000000111000000",
		10 => "000000111000000111000000",
		11 => "000000111000000111000000",
		12 => "000000111000000111000000",
		13 => "000000011100001110000000",
		14 => "000000001111111100000000",
		15 => "000000000111111000000000",
		16 => "000000011111111110000000",
		17 => "000000111100001111000000",
		18 => "000000111000000111000000",
		19 => "000001110000000011100000",
		20 => "000001110000000011100000",
		21 => "000001110000000011100000",
		22 => "000001111000000111100000",
		23 => "000001111100001111000000",
		24 => "000000111111111111000000",
		25 => "000000011111111110000000",
		26 => "000000000111111000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	constant rom_mdl_9 : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000001111110000000000",
		 6 => "000000111111111000000000",
		 7 => "000001111111111100000000",
		 8 => "000001111000011110000000",
		 9 => "000011110000001110000000",
		10 => "000011100000000110000000",
		11 => "000011100000000111000000",
		12 => "000011100000000111000000",
		13 => "000011100000000111000000",
		14 => "000011110000001111000000",
		15 => "000001111000011111000000",
		16 => "000001111111110111000000",
		17 => "000000111111110111000000",
		18 => "000000001111000111000000",
		19 => "000000000000000111000000",
		20 => "000000000000001111000000",
		21 => "000000000000001110000000",
		22 => "000000000000011110000000",
		23 => "000000100000111100000000",
		24 => "000000111111111100000000",
		25 => "000000111111111000000000",
		26 => "000000011111100000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
	
	constant rom_mdl_dp : rom_mem_t := (
		 0 => "000000000000000000000000",
		 1 => "000000000000000000000000",
		 2 => "000000000000000000000000",
		 3 => "000000000000000000000000",
		 4 => "000000000000000000000000",
		 5 => "000000000000000000000000",
		 6 => "000000000000000000000000",
		 7 => "000000000000000000000000",
		 8 => "000000000000000000000000",
		 9 => "000000000001100000000000",
		10 => "000000000011110000000000",
		11 => "000000000011110000000000",
		12 => "000000000001100000000000",
		13 => "000000000000000000000000",
		14 => "000000000000000000000000",
		15 => "000000000000000000000000",
		16 => "000000000000000000000000",
		17 => "000000000000000000000000",
		18 => "000000000000000000000000",
		19 => "000000000000000000000000",
		20 => "000000000001100000000000",
		21 => "000000000011110000000000",
		22 => "000000000011110000000000",
		23 => "000000000001100000000000",
		24 => "000000000000000000000000",
		25 => "000000000000000000000000",
		26 => "000000000000000000000000",
		27 => "000000000000000000000000",
		28 => "000000000000000000000000",
		29 => "000000000000000000000000",
		30 => "000000000000000000000000",
		31 => "000000000000000000000000");
		
	signal bit_dat	: std_logic_vector(0 to ROM_WIDTH - 1);
	signal num_adr	: std_logic_vector(3 downto 0);
	signal bit_adr	: std_logic_vector(4 downto 0);
	
begin
	
	num_adr <= rom_adr_i(8 downto 5);
	bit_adr <= rom_adr_i(4 downto 0);
	
	process(num_adr, bit_adr, bit_dat)
	begin
		case num_adr is
			when "0000" => bit_dat <= rom_mdl_0(to_integer(unsigned(bit_adr)));
			when "0001" => bit_dat <= rom_mdl_1(to_integer(unsigned(bit_adr)));
			when "0010" => bit_dat <= rom_mdl_2(to_integer(unsigned(bit_adr)));
			when "0011" => bit_dat <= rom_mdl_3(to_integer(unsigned(bit_adr)));
			when "0100" => bit_dat <= rom_mdl_4(to_integer(unsigned(bit_adr)));
			when "0101" => bit_dat <= rom_mdl_5(to_integer(unsigned(bit_adr)));
			when "0110" => bit_dat <= rom_mdl_6(to_integer(unsigned(bit_adr)));
			when "0111" => bit_dat <= rom_mdl_7(to_integer(unsigned(bit_adr)));
			when "1000" => bit_dat <= rom_mdl_8(to_integer(unsigned(bit_adr)));
			when "1001" => bit_dat <= rom_mdl_9(to_integer(unsigned(bit_adr)));
			when "1010" => bit_dat <= rom_mdl_dp(to_integer(unsigned(bit_adr)));
			when others => bit_dat <= (others => '0');
		end case;
		
		rom_dat_o <= bit_dat;
	end process;
end rtl;